
/****************************************************************************
 * fwperiph_dma.sv
 ****************************************************************************/

  
/**
 * Module: fwperiph_dma
 * 
 * TODO: Add module documentation
 */
module fwperiph_dma #(
		);


endmodule


