/****************************************************************************
 * sv_bfms_api_pkg.sv
 ****************************************************************************/

/**
 * Package: sv_bfms_api_pkg
 * 
 * TODO: Add package documentation
 */
package sv_bfms_api_pkg;
	`include "sv_bfms_rw_api_if.svh"

endpackage


