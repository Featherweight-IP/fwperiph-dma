/****************************************************************************
 * wb_dma_coverage_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: wb_dma_coverage_pkg
 * 
 * TODO: Add package documentation
 */
package wb_dma_coverage_pkg;
	import uvm_pkg::*;
	import wb_dma_env_pkg::*;

	`include "wb_dma_single_transfer_descriptor_cov.svh"

endpackage


