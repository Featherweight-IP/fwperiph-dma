/****************************************************************************
 * wb_dma_ll_transfer_descriptor.svh
 ****************************************************************************/

/**
 * Class: wb_dma_ll_transfer_descriptor
 * 
 * TODO: Add class documentation
 */
class wb_dma_ll_transfer_descriptor extends wb_dma_descriptor;
	`uvm_object_utils(wb_dma_ll_transfer_descriptor)

//	// disable linked-list transfers
//	constraint ll_desc_sz_c {
//		ll_desc_sz == 4;
//	}
//	
//	constraint transfer_sz_c {
//		transfer_sz == 16;
//	}

endclass


