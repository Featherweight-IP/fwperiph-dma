/****************************************************************************
 *  mem_mgr_pkg.sv
 ****************************************************************************/

`include "uvm_macros.svh"
package mem_mgr_pkg;
	import uvm_pkg::*;
	`include "mem_mgr_ev.svh"
	`include "mem_mgr.svh"
endpackage
