
/****************************************************************************
 * fwperiph_dma_dbg.v
 ****************************************************************************/

  
/**
 * Module: fwperiph_dma_dbg
 * 
 * TODO: Add module documentation
 */
module fwperiph_dma_dbg #(
		parameter ch_count=1
		) (
		input				clock,
		input[31:0]			adr,
		input[31:0]			dat_w,
		input[31:0]			we
		);

	// Empty

endmodule


