
/****************************************************************************
 * fwperiph_dma_wb_4.v
 ****************************************************************************/

  
/**
 * Module: fwperiph_dma_wb_4
 * 
 * TODO: Add module documentation
 */
module fwperiph_dma_wb_4;


endmodule


